`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.04.2024 15:07:20
// Design Name: 
// Module Name: cla_16bit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module cla_16bit(A, B, Cin, S, Cout);
input [15:0]A, B;
input Cin;
output [15:0] S;
output Cout;

  wire P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15;
  wire [15:0] Ci;
  
  // P Stage
  assign P0 = A[0] ^ B[0];
  assign P1 = A[1] ^ B[1];
  assign P2 = A[2] ^ B[2];
  assign P3 = A[3] ^ B[3];
  assign P4 = A[4] ^ B[4];
  assign P5 = A[5] ^ B[5];
  assign P6 = A[6] ^ B[6];
  assign P7 = A[7] ^ B[7];
  assign P8 = A[8] ^ B[8];
  assign P9 = A[9] ^ B[9];
  assign P10 = A[10] ^ B[10];
  assign P11 = A[11] ^ B[11];
  assign P12 = A[12] ^ B[12];
  assign P13 = A[13] ^ B[13];
  assign P14 = A[14] ^ B[14];
  assign P15 = A[15] ^ B[15];
 
  //Carry Stage
  assign Ci[0] = Cin;
  assign Ci[1] = (A[0] & B[0]) | ((A[0]^B[0]) & Ci[0]);
  assign Ci[2] = (A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])));
  assign Ci[3] = (A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))));
  assign Ci[4] = (A[3] & B[3]) | ((A[3]^B[3]) & ((A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))))));
  assign Ci[5] = (A[4] & B[4]) | ((A[4]^B[4]) & ((A[3] & B[3]) | ((A[3]^B[3]) & ((A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))))))));
  assign Ci[6] = (A[5] & B[5]) | ((A[5]^B[5]) & ((A[4] & B[4]) | ((A[4]^B[4]) & ((A[3] & B[3]) | ((A[3]^B[3]) & ((A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))))))))));
  assign Ci[7] = (A[6] & B[6]) | ((A[6]^B[6]) & ((A[5] & B[5]) | ((A[5]^B[5]) & ((A[4] & B[4]) | ((A[4]^B[4]) & ((A[3] & B[3]) | ((A[3]^B[3]) & ((A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))))))))))));
  assign Ci[8] = (A[7] & B[7]) | ((A[7]^B[7]) & ((A[6] & B[6]) | ((A[6]^B[6]) & ((A[5] & B[5]) | ((A[5]^B[5]) & ((A[4] & B[4]) | ((A[4]^B[4]) & ((A[3] & B[3]) | ((A[3]^B[3]) & ((A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))))))))))))));
  assign Ci[9] = (A[8] & B[8]) | ((A[8]^B[8]) & ((A[7] & B[7]) | ((A[7]^B[7]) & ((A[6] & B[6]) | ((A[6]^B[6]) & ((A[5] & B[5]) | ((A[5]^B[5]) & ((A[4] & B[4]) | ((A[4]^B[4]) & ((A[3] & B[3]) | ((A[3]^B[3]) & ((A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))))))))))))))));
  assign Ci[10] = (A[9] & B[9]) | ((A[9]^B[9]) & ((A[8] & B[8]) | ((A[8]^B[8]) & ((A[7] & B[7]) | ((A[7]^B[7]) & ((A[6] & B[6]) | ((A[6]^B[6]) & ((A[5] & B[5]) | ((A[5]^B[5]) & ((A[4] & B[4]) | ((A[4]^B[4]) & ((A[3] & B[3]) | ((A[3]^B[3]) & ((A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))))))))))))))))));
  assign Ci[11] = (A[10] & B[10]) | ((A[10]^B[10]) & ((A[9] & B[9]) | ((A[9]^B[9]) & ((A[8] & B[8]) | ((A[8]^B[8]) & ((A[7] & B[7]) | ((A[7]^B[7]) & ((A[6] & B[6]) | ((A[6]^B[6]) & ((A[5] & B[5]) | ((A[5]^B[5]) & ((A[4] & B[4]) | ((A[4]^B[4]) & ((A[3] & B[3]) | ((A[3]^B[3]) & ((A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))))))))))))))))))));
  assign Ci[12] = (A[11] & B[11]) | ((A[11]^B[11]) & ((A[10] & B[10]) | ((A[10]^B[10]) & ((A[9] & B[9]) | ((A[9]^B[9]) & ((A[8] & B[8]) | ((A[8]^B[8]) & ((A[7] & B[7]) | ((A[7]^B[7]) & ((A[6] & B[6]) | ((A[6]^B[6]) & ((A[5] & B[5]) | ((A[5]^B[5]) & ((A[4] & B[4]) | ((A[4]^B[4]) & ((A[3] & B[3]) | ((A[3]^B[3]) & ((A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))))))))))))))))))))));
  assign Ci[13] = (A[12] & B[12]) | ((A[12]^B[12]) & ((A[11] & B[11]) | ((A[11]^B[11]) & ((A[10] & B[10]) | ((A[10]^B[10]) & ((A[9] & B[9]) | ((A[9]^B[9]) & ((A[8] & B[8]) | ((A[8]^B[8]) & ((A[7] & B[7]) | ((A[7]^B[7]) & ((A[6] & B[6]) | ((A[6]^B[6]) & ((A[5] & B[5]) | ((A[5]^B[5]) & ((A[4] & B[4]) | ((A[4]^B[4]) & ((A[3] & B[3]) | ((A[3]^B[3]) & ((A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))))))))))))))))))))))));
  assign Ci[14] = (A[13] & B[13]) | ((A[13]^B[13]) & ((A[12] & B[12]) | ((A[12]^B[12]) & ((A[11] & B[11]) | ((A[11]^B[11]) & ((A[10] & B[10]) | ((A[10]^B[10]) & ((A[9] & B[9]) | ((A[9]^B[9]) & ((A[8] & B[8]) | ((A[8]^B[8]) & ((A[7] & B[7]) | ((A[7]^B[7]) & ((A[6] & B[6]) | ((A[6]^B[6]) & ((A[5] & B[5]) | ((A[5]^B[5]) & ((A[4] & B[4]) | ((A[4]^B[4]) & ((A[3] & B[3]) | ((A[3]^B[3]) & ((A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))))))))))))))))))))))))));
  assign Ci[15] = (A[14] & B[14]) | ((A[14]^B[14]) & ((A[13] & B[13]) | ((A[13]^B[13]) & ((A[12] & B[12]) | ((A[12]^B[12]) & ((A[11] & B[11]) | ((A[11]^B[11]) & ((A[10] & B[10]) | ((A[10]^B[10]) & ((A[9] & B[9]) | ((A[9]^B[9]) & ((A[8] & B[8]) | ((A[8]^B[8]) & ((A[7] & B[7]) | ((A[7]^B[7]) & ((A[6] & B[6]) | ((A[6]^B[6]) & ((A[5] & B[5]) | ((A[5]^B[5]) & ((A[4] & B[4]) | ((A[4]^B[4]) & ((A[3] & B[3]) | ((A[3]^B[3]) & ((A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))))))))))))))))))))))))))));
  assign Cout  = (A[15] & B[15]) | ((A[15]^B[15]) & ((A[14] & B[14]) | ((A[14]^B[14]) & ((A[13] & B[13]) | ((A[13]^B[13]) & ((A[12] & B[12]) | ((A[12]^B[12]) & ((A[11] & B[11]) | ((A[11]^B[11]) & ((A[10] & B[10]) | ((A[10]^B[10]) & ((A[9] & B[9]) | ((A[9]^B[9]) & ((A[8] & B[8]) | ((A[8]^B[8]) & ((A[7] & B[7]) | ((A[7]^B[7]) & ((A[6] & B[6]) | ((A[6]^B[6]) & ((A[5] & B[5]) | ((A[5]^B[5]) & ((A[4] & B[4]) | ((A[4]^B[4]) & ((A[3] & B[3]) | ((A[3]^B[3]) & ((A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))))))))))))))))))))))))))))));
  
  // Sum Stage
  assign S[0] = P0 ^ Cin;
  assign S[1] = P1 ^ Ci[1];
  assign S[2] = P2 ^ Ci[2];
  assign S[3] = P3 ^ Ci[3];
  assign S[4] = P4 ^ Ci[4]; 
  assign S[5] = P5 ^ Ci[5];
  assign S[6] = P6 ^ Ci[6];
  assign S[7] = P7 ^ Ci[7];
  assign S[8] = P8 ^ Ci[8];
  assign S[9] = P9 ^ Ci[9];
  assign S[10] = P10 ^ Ci[10];
  assign S[11] = P11 ^ Ci[11];
  assign S[12] = P12 ^ Ci[12];
  assign S[13] = P13 ^ Ci[13];
  assign S[14] = P14 ^ Ci[14];
  assign S[15] = P15 ^ Ci[15];
  
endmodule
